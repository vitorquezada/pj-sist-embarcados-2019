module detectorDeCancer(IO, reset, HEX5, HEX3, HEX2, HEX1, HEX0);

	
    
endmodule
